// issp.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module issp (
		output wire [1:0] source  // sources.source
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("INIT"),
		.probe_width             (0),
		.source_width            (2),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (source), // sources.source
		.source_ena (1'b1)    // (terminated)
	);

endmodule
