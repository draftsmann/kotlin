
module rst_button (
	source);	

	output	[0:0]	source;
endmodule
