
module issp_sel_data (
	source);	

	output	[0:0]	source;
endmodule
