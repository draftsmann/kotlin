
module issp (
	source);	

	output	[1:0]	source;
endmodule
